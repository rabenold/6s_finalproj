`timescale 1ns / 1ps
`default_nettype none
    module zig_zagger #(parameter DATA_WIDTH = 11, WITDH = 8, HEIGHT = 8)(
        input logic [DATA_WIDTH-1:0] input_matrix [0:WIDTH-1][0:HEIGHT-1],
        output logic [DATA_WIDTH-1:0] zig_zag_out [63:0],
    )
    //define the first element as 0 using this notation 

 always_comb begin
        // For each zig-zag index, directly assign the corresponding matrix value
        zig_zag_out[0]  = input_matrix[0][0];  // (0,0)
        zig_zag_out[1]  = input_matrix[0][1];  // (0,1)
        zig_zag_out[2]  = input_matrix[1][0];  // (1,0)
        zig_zag_out[3]  = input_matrix[2][0];  // (2,0)
        zig_zag_out[4]  = input_matrix[1][1];  // (1,1)
        zig_zag_out[5]  = input_matrix[0][2];  // (0,2)
        zig_zag_out[6]  = input_matrix[0][3];  // (0,3)
        zig_zag_out[7]  = input_matrix[1][2];  // (1,2)
        zig_zag_out[8]  = input_matrix[2][1];  // (2,1)
        zig_zag_out[9]  = input_matrix[3][0];  // (3,0)
        zig_zag_out[10] = input_matrix[4][0];  // (4,0)
        zig_zag_out[11] = input_matrix[3][1];  // (3,1)
        zig_zag_out[12] = input_matrix[2][2];  // (2,2)
        zig_zag_out[13] = input_matrix[1][3];  // (1,3)
        zig_zag_out[14] = input_matrix[0][4];  // (0,4)
        zig_zag_out[15] = input_matrix[0][5];  // (0,5)
        zig_zag_out[16] = input_matrix[1][4];  // (1,4)
        zig_zag_out[17] = input_matrix[2][3];  // (2,3)
        zig_zag_out[18] = input_matrix[3][2];  // (3,2)
        zig_zag_out[19] = input_matrix[4][1];  // (4,1)
        zig_zag_out[20] = input_matrix[5][0];  // (5,0)
        zig_zag_out[21] = input_matrix[6][0];  // (6,0)
        zig_zag_out[22] = input_matrix[5][1];  // (5,1)
        zig_zag_out[23] = input_matrix[4][2];  // (4,2)
        zig_zag_out[24] = input_matrix[3][3];  // (3,3)
        zig_zag_out[25] = input_matrix[2][4];  // (2,4)
        zig_zag_out[26] = input_matrix[1][5];  // (1,5)
        zig_zag_out[27] = input_matrix[0][6];  // (0,6)
        zig_zag_out[28] = input_matrix[0][7];  // (0,7)
        zig_zag_out[29] = input_matrix[1][6];  // (1,6)
        zig_zag_out[30] = input_matrix[2][5];  // (2,5)
        zig_zag_out[31] = input_matrix[3][4];  // (3,4)
        zig_zag_out[32] = input_matrix[4][3];  // (4,3)
        zig_zag_out[33] = input_matrix[5][2];  // (5,2)
        zig_zag_out[34] = input_matrix[6][1];  // (6,1)
        zig_zag_out[35] = input_matrix[7][0];  // (7,0)
        zig_zag_out[36] = input_matrix[7][1];  // (7,1)
        zig_zag_out[37] = input_matrix[6][2];  // (6,2)
        zig_zag_out[38] = input_matrix[5][3];  // (5,3)
        zig_zag_out[39] = input_matrix[4][4];  // (4,4)
        zig_zag_out[40] = input_matrix[3][5];  // (3,5)
        zig_zag_out[41] = input_matrix[2][6];  // (2,6)
        zig_zag_out[42] = input_matrix[1][7];  // (1,7)
        zig_zag_out[43] = input_matrix[2][7];  // (2,7)
        zig_zag_out[44] = input_matrix[3][6];  // (3,6)
        zig_zag_out[45] = input_matrix[4][5];  // (4,5)
        zig_zag_out[46] = input_matrix[5][4];  // (5,4)
        zig_zag_out[47] = input_matrix[6][3];  // (6,3)
        zig_zag_out[48] = input_matrix[7][2];  // (7,2)
        zig_zag_out[49] = input_matrix[7][3];  // (7,3)
        zig_zag_out[50] = input_matrix[6][4];  // (6,4)
        zig_zag_out[51] = input_matrix[5][5];  // (5,5)
        zig_zag_out[52] = input_matrix[4][6];  // (4,6)
        zig_zag_out[53] = input_matrix[3][7];  // (3,7)
        zig_zag_out[54] = input_matrix[4][7];  // (4,7)
        zig_zag_out[55] = input_matrix[5][6];  // (5,6)
        zig_zag_out[56] = input_matrix[6][5];  // (6,5)
        zig_zag_out[57] = input_matrix[7][4];  // (7,4)
        zig_zag_out[58] = input_matrix[7][5];  // (7,5)
        zig_zag_out[59] = input_matrix[6][6];  // (6,6)
        zig_zag_out[60] = input_matrix[5][7];  // (5,7)
        zig_zag_out[61] = input_matrix[6][7];  // (6,7)
        zig_zag_out[62] = input_matrix[7][6];  // (7,6)
        zig_zag_out[63] = input_matrix[7][7];  // (7,7)
    end
endmodule
`default_nettype wire

