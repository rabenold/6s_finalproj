`timescale 1ns / 1ps
`default_nettype none





`default_nettype wire // prevents system from inferring an undeclared logic (good practice)
