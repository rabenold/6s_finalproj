`timescale 1ns / 1ps
`default_nettype none
    module buffer_slicer #(parameter DATA_WIDTH = 16)(
    input logic [8:0] x_in,
    input logic [8:0] y_in    

    output [DATA_WIDTH-1:0] logic [DATA_WIDTH-1:0] matrix_out
 
    )
     
     
    endmodule

`default_nettype wire

